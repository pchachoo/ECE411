--
-- VHDL Architecture ece411.DRAM.untitled
--
-- Created:
--          by - chachon2.ews (linux-a1.ews.illinois.edu)
--          at - 20:36:55 08/02/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY DRAM IS
-- Declarations

END DRAM ;

--
ARCHITECTURE untitled OF DRAM IS
BEGIN
END ARCHITECTURE untitled;

